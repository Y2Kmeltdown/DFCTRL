module spi_top #(
    parameter 
    WIDTH_ADDR_ACT = 11, 
    WIDTH_ACT_MEM = 8, 
    ACT_MEM_HEADER = 8'b10,
    
    WIDTH_ADDR_PARAM = 13, 
    WIDTH_PARAM_MEM = 128,
    PARAM_MEM_HEADER = 8'b01,

    WIDTH_ADDR_INST = 6,
    WIDTH_INST_MEM = 80, 
    INST_MEM_HEADER = 8'b11,
     
    WIDTH_SPI_WORD = 8,
    SPI_OUT_ADDRESS_SIZE = 4,
    SPI_IN_ADDRESS_SIZE = 4,
    SPI_OUT_ADDRESS_DEPTH = 16
) 
(
    input   reset_n,
    input   clk,


    input   spi_clk,
    input   MOSI,
    output  MISO,
    input   chip_select_n,
    input   [1:0]   set_reg,

    output  [WIDTH_ADDR_ACT-1:0]    act_mem_addr,
    output  [WIDTH_ACT_MEM-1:0]     act_mem_data,
    output                          act_mem_wren,
    input   [WIDTH_ACT_MEM-1:0]     act_mem_q,
    output                          data_ready,
    output                          sel_ext,

    output  [WIDTH_ADDR_PARAM-1:0]  param_mem_addr,
    output  [WIDTH_PARAM_MEM-1:0]   param_mem_data,
    output                          param_mem_wren,

    output  [WIDTH_ADDR_INST-1:0]   inst_mem_addr,
    output  [WIDTH_INST_MEM-1:0]    inst_mem_data,
    output                          inst_mem_wren,

    output                          proc_enable,
    output                          proc_reset

    // Inputs data from system
);

wire [7:0]  internal_in;
wire        wr_req;
wire        write_full;
wire        write_empty;


wire [7:0]  internal_out;
wire        rd_req;
wire        read_full;
wire        read_empty;


spi_controller #(
    .SPI_BUS_WIDTH(WIDTH_SPI_WORD),
    .SPI_OUT_ADDRESS_SIZE(SPI_OUT_ADDRESS_SIZE),
    .SPI_IN_ADDRESS_SIZE(SPI_IN_ADDRESS_SIZE)
) 
    spi_controller_0 (
    .reset_n(reset_n),

    .spi_clk(spi_clk),
    .mosi(MOSI),
    .miso(MISO),
    .chip_select_n(chip_select_n),
    .set_reg(set_reg),
    
    .wr_req(wr_req),
    .internal_clk(clk),
    .internal_in(act_mem_q),
    .SPI_write_full(write_full),
    .SPI_write_empty(write_empty),

    .internal_out(internal_out),
    .rd_req(rd_req),
    .SPI_read_full(read_full),
    .SPI_read_empty(read_empty)
);

packetizer #(
    .WIDTH_ADDR_ACT(WIDTH_ADDR_ACT), 
    .WIDTH_ACT_MEM(WIDTH_ACT_MEM), 
    .ACT_MEM_HEADER(ACT_MEM_HEADER),
    
    .WIDTH_ADDR_PARAM(WIDTH_ADDR_PARAM), 
    .WIDTH_PARAM_MEM(WIDTH_PARAM_MEM),
    .PARAM_MEM_HEADER(PARAM_MEM_HEADER),

    .WIDTH_ADDR_INST(WIDTH_ADDR_INST),
    .WIDTH_INST_MEM(WIDTH_INST_MEM), 
    .INST_MEM_HEADER(INST_MEM_HEADER),
     
    .WIDTH_SPI_WORD(WIDTH_SPI_WORD),
    .SPI_OUT_ADDRESS_SIZE(SPI_OUT_ADDRESS_SIZE),
    .SPI_IN_ADDRESS_SIZE(SPI_IN_ADDRESS_SIZE),
    .SPI_OUT_ADDRESS_DEPTH(SPI_OUT_ADDRESS_DEPTH)
)
packetizer_0
(
    .reset_n(reset_n),
    .clk(clk),
    .spi_clk(spi_clk),
    .chip_select_n(chip_select_n),

    .spi_word(internal_out),
    .read_fifo_empty(read_empty),
    .write_fifo_empty(write_empty),
    .write_fifo_full(write_full),
    .rd_req(rd_req),
    .wr_req(wr_req),
    .sel_ext(sel_ext),

    .act_mem_addr(act_mem_addr),
    .act_mem_data(act_mem_data),
    .act_mem_wren(act_mem_wren),
    .data_ready(data_ready),


    .param_mem_addr(param_mem_addr),
    .param_mem_data(param_mem_data),
    .param_mem_wren(param_mem_wren),

    .inst_mem_addr(inst_mem_addr),
    .inst_mem_data(inst_mem_data),
    .inst_mem_wren(inst_mem_wren),

    .proc_enable(proc_enable),
    .proc_reset(proc_reset)
);

// Module for writing to SPI bus


endmodule